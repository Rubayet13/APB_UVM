package env_pkg;

  import agent_pkg::*;
  
  `include "../tb_top/params.sv"
  `include "apb_sco.sv"
  `include "apb_env.sv"

endpackage