package agent_pkg;

    `include "../tb/tb_top/params.sv"
    `include "apb_trans.sv"
    `include "apb_config.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_agent.sv"

endpackage